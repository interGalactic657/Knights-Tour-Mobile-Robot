/////////////////////////////////////////////////
// inert_intf_tb.sv                           //
// This testbench simulates calibrating the  //
// the 6-axis DEO Nano gyro.                //
/////////////////////////////////////////////
module inert_intf_tb();

  logic clk, rst_n; // Clock and reset signals.
  logic SS_n; // Active low chip select for SPI communication.
  logic strt_cal, cal_done; // Signals to start and indicate completion of calibration.
  logic SCLK, MOSI, MISO; // SPI clock, MOSI (Master Out Serf In), and MISO (Master In Serf Out) signals.
  logic INT; // Interrupt signal from the inertial sensor.
  logic rdy; // Ready signal indicating sensor is ready for measurement.
  logic [11:0] heading; // 12-bit heading value from the sensor.

  //////////////////////////////////////////
  // Instantiate the inertal system DUTs //
  ////////////////////////////////////////
  // Instantiate the inertial interface (iINERT) module.
  inert_intf iINERT(
    .clk(clk), .rst_n(rst_n), .strt_cal(strt_cal), .cal_done(cal_done), 
    .heading(heading), .rdy(rdy), .lftIR(1'b0), .rghtIR(1'b0), 
    .SS_n(SS_n), .SCLK(SCLK), .MOSI(MOSI), .MISO(MISO), .INT(INT),
    .moving(1'b1)
  );

  // Instantiate the NEMO gyro sensor (iNEMO).
  SPI_iNEMO2 iNEMO(
    .SS_n(SS_n), .SCLK(SCLK), .MISO(MISO), .MOSI(MOSI), .INT(INT)
  );
  /////////////////////////////////////////////////////////////////////

  ////////////////////////////////////////////////////////////
  // Task to wait for a signal to be asserted, otherwise   //
  // times out.                                           //
  /////////////////////////////////////////////////////////
  task automatic timeout_task(ref sig, input int clks2wait, input string signal);
    fork
      begin : timeout
        repeat(clks2wait) @(posedge clk);
        $display("ERROR: %s not getting asserted and/or held at its value.", signal);
        $stop(); // Stop simulation on error.
      end : timeout
      begin
        @(posedge sig) disable timeout; // Disable timeout if sig is asserted.
      end
    join
  endtask

  ///////////////////////////////////////////////////////////
  // Apply stimulus and check response as to whether an    //
  // interrupt is being generated by the inertial          //
  // sensor as well as whether calibration was successful. //
  ///////////////////////////////////////////////////////////
  initial begin
    clk = 1'b0; // initially clock is low
		rst_n = 1'b0; // reset the system
    strt_cal = 1'b0; // Do not start calibration initially.
    
     // Wait 1.5 clocks for reset
    @(posedge clk);
    @(negedge clk) rst_n = 1'b1; // Deassert reset on a negative edge of clock

    ///////////////////////////////////////////////////////
    // TEST 1: Check that NEMO's setup signal goes high //
    /////////////////////////////////////////////////////
    // Wait for NEMO_setup to be asserted, or timeout after a 100000 clocks.
    fork
      begin : timeout_setup
        repeat(1000000) @(posedge clk);
        $display("ERROR: NEMO_setup not getting asserted and/or held at its value.");
        $stop(); // Stop simulation on error.
      end : timeout_setup
      begin
        @(posedge iNEMO.NEMO_setup) disable timeout_setup; // Disable timeout if NEMO_setup is asserted.
      end
    join

    /////////////////////////////////////////////////////
    // TEST 2: Check that cal_done signal is asserted //
    ///////////////////////////////////////////////////
    // Start calibration process by asserting strt_cal.
    @(negedge clk) strt_cal = 1'b1; // Begin calibration on negative edge of clock.
    @(negedge clk) strt_cal = 1'b0; // Deassert strt_cal after one clock.

    // Wait for cal_done to be asserted, or timeout after a 1000000 clocks.
    timeout_task(.sig(cal_done), .clks2wait(1000000), .signal("cal_done"));

    // Let the simulation run for an additional 8 million clock cycles to generate waveforms.
    repeat(8000000) @(posedge clk);

    // End the simulation after waveform generation.
    $stop();
  end

  always
    #5 clk = ~clk; // toggle clock every 5 time units
endmodule
